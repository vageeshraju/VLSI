module half_subtractor(output d,bor, input a,b);
assign d = a^b;
assign bor= (~a) & b;
endmodule
