module full_adder_tb();
reg a,b,cin;
wire sum,carry;
full_adder dut (
.a(a),
.b(b),
.cin(cin),
.sum(sum),
.carry(carry));
initial begin
$dumpfile ("fulladder.vcd");
$dumpvars (0,full_adder_tb);
  $monitor ("a=%b,b=%b,cin=%b,sum=%b,carry=%b",a,b,cin,sum,carry);
#5a=0;b=0;cin=0;
#5a=0;b=1;cin=0;
#5a=1;b=0;cin=0;
#5a=1;b=1;cin=0;
#5a=0;b=0;cin=1;
#5a=0;b=1;cin=1;
#5a=1;b=0;cin=1;
#5a=1;b=1;cin=1;
#40 $finish;
end
endmodule
