module not (
    output y,
    input a
);
assign y=~a;
endmodule
