`timescale 1ns/1ps
module encoder8X3_tb();
 wire x1,x2,x3;
 reg i0,i1,i2,i3,i4,i5,i6,i7;
encoder8X3 dut (
.x1(x1),
.x2(x2),
.x3(x3),
.i0(i0),
.i1(i1),
.i2(i2),
.i3(i3),
.i4(i4),
.i5(i5),
.i6(i6),
.i7(i7));
initial begin
$dumpfile("encoder8X3.vcd");
$dumpvars (0,encoder8X3_tb);
$monitor ("time=%t,x3=%b,x2=%b,x1=%b,i0=%b,i1=%b,i2=%b,i3=%b,i4=%b,i5=%b,i6=%b,i7=%b",$time,x3,x2,x1,i0,i1,i2,i3,i4,i5,i6,i7);
#5i0=1;i1=0;i2=0;i3=0;i4=0;i5=0;i6=0;i7=0;
#5i0=0;i1=1;i2=0;i3=0;i4=0;i5=0;i6=0;i7=0;
#5i0=0;i1=0;i2=1;i3=0;i4=0;i5=0;i6=0;i7=0;
#5i0=0;i1=0;i2=0;i3=1;i4=0;i5=0;i6=0;i7=0;
#5i0=0;i1=0;i2=0;i3=0;i4=1;i5=0;i6=0;i7=0;
#5i0=0;i1=0;i2=0;i3=0;i4=0;i5=1;i6=0;i7=0;
#5i0=0;i1=0;i2=0;i3=0;i4=0;i5=0;i6=1;i7=0;
#5i0=0;i1=0;i2=0;i3=0;i4=0;i5=0;i6=0;i7=1;
#40$finish;
end
endmodule
