module exor_gate (
    output x,
    input a,b
);
assign x=a^b;
endmodule
